* Simple resistor divider
V1 1 0 DC 10
R1 1 2 1k
R2 2 0 2k
.end
